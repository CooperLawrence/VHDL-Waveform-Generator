library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity Memory is
port(
	CS: in std_logic_vector(1 downto 0); --Current state
	EN: in std_logic; --Enable
	dataBus: out std_logic_vector(31 downto 0); --Data Bus
	address: in std_logic_vector (6 downto 0) -- Address bus
	);
end Memory;

architecture MemArch of Memory is
type Sine_array is array (0 to 127) of integer; --look-up table for Sine wave
type Square_array is array (0 to 127) of integer; --look-up table for Square wave
type Triangle_array is array (0 to 127) of integer; --look-up table for Triangle wave
type Special_array is array (0 to 127) of integer; --look-up table for damped-sine wave

signal sine : Sine_array;
signal square : Square_array;
signal triangle : Triangle_array;
signal special : Special_array;



begin
sine <= (0 ,
6 ,
12 ,
18 ,
24 ,
31 ,
37 ,
43 ,
48 ,
54 ,
60 ,
65 ,
71 ,
76 ,
81 ,
85 ,
90 ,
94 ,
98 ,
102 ,
106 ,
109 ,
112 ,
115 ,
118 ,
120 ,
122 ,
124 ,
125 ,
126 ,
127 ,
127 ,
128 ,
127 ,
127 ,
126 ,
125 ,
124 ,
122 ,
120 ,
118 ,
115 ,
112 ,
109 ,
106 ,
102 ,
98 ,
94 ,
90 ,
85 ,
81 ,
76 ,
71 ,
65 ,
60 ,
54 ,
48 ,
43 ,
37 ,
31 ,
24 ,
18 ,
12 ,
6 ,
0 ,
-6 ,
-12 ,
-18 ,
-24 ,
-31 ,
-37 ,
-43 ,
-48 ,
-54 ,
-60 ,
-65 ,
-71 ,
-76 ,
-81 ,
-85 ,
-90 ,
-94 ,
-98 ,
-102 ,
-106 ,
-109 ,
-112 ,
-115 ,
-118 ,
-120 ,
-122 ,
-124 ,
-125 ,
-126 ,
-127 ,
-127 ,
-128 ,
-127 ,
-127 ,
-126 ,
-125 ,
-124 ,
-122 ,
-120 ,
-118 ,
-115 ,
-112 ,
-109 ,
-106 ,
-102 ,
-98 ,
-94 ,
-90 ,
-85 ,
-81 ,
-76 ,
-71 ,
-65 ,
-60 ,
-54 ,
-48 ,
-43 ,
-37 ,
-31 ,
-24 ,
-18 ,
-12 ,
-6);
square <= (128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128 ,
-128);
triangle <= (0 ,
4 ,
8 ,
12 ,
16 ,
20 ,
24 ,
28 ,
32 ,
36 ,
40 ,
44 ,
48 ,
52 ,
56 ,
60 ,
64 ,
68 ,
72 ,
76 ,
80 ,
84 ,
88 ,
92 ,
96 ,
100 ,
104 ,
108 ,
112 ,
116 ,
120 ,
124 ,
128 ,
124 ,
120 ,
116 ,
112 ,
108 ,
104 ,
100 ,
96 ,
92 ,
88 ,
84 ,
80 ,
76 ,
72 ,
68 ,
64 ,
60 ,
56 ,
52 ,
48 ,
44 ,
40 ,
36 ,
32 ,
28 ,
24 ,
20 ,
16 ,
12 ,
8 ,
4 ,
0 ,
-4 ,
-8 ,
-12 ,
-16 ,
-20 ,
-24 ,
-28 ,
-32 ,
-36 ,
-40 ,
-44 ,
-48 ,
-52 ,
-56 ,
-60 ,
-64 ,
-68 ,
-72 ,
-76 ,
-80 ,
-84 ,
-88 ,
-92 ,
-96 ,
-100 ,
-104 ,
-108 ,
-112 ,
-116 ,
-120 ,
-124 ,
0 ,
4 ,
8 ,
12 ,
16 ,
20 ,
24 ,
28 ,
32 ,
36 ,
40 ,
44 ,
48 ,
52 ,
56 ,
60 ,
64 ,
68 ,
72 ,
76 ,
80 ,
84 ,
88 ,
92 ,
96 ,
100 ,
104 ,
108 ,
112 ,
116 ,
120 ,
124);
special <= (0 ,
0 ,
0 ,
0 ,
0 ,
1 ,
1 ,
2 ,
3 ,
3 ,
4 ,
5 ,
6 ,
7 ,
8 ,
10 ,
11 ,
12 ,
13 ,
15 ,
16 ,
18 ,
19 ,
20 ,
22 ,
23 ,
24 ,
26 ,
27 ,
28 ,
29 ,
30 ,
32 ,
32 ,
33 ,
34 ,
35 ,
35 ,
36 ,
36 ,
36 ,
37 ,
37 ,
36 ,
36 ,
36 ,
35 ,
34 ,
33 ,
32 ,
31 ,
30 ,
28 ,
27 ,
25 ,
23 ,
21 ,
19 ,
16 ,
14 ,
11 ,
8 ,
6 ,
3 ,
0 ,
-3 ,
-6 ,
-9 ,
-13 ,
-16 ,
-20 ,
-23 ,
-27 ,
-31 ,
-34 ,
-38 ,
-42 ,
-45 ,
-49 ,
-53 ,
-56 ,
-60 ,
-63 ,
-66 ,
-69 ,
-72 ,
-75 ,
-78 ,
-81 ,
-83 ,
-86 ,
-88 ,
-90 ,
-91 ,
-93 ,
-94 ,
-96 ,
-96 ,
-97 ,
-97 ,
-98 ,
-97 ,
-97 ,
-96 ,
-96 ,
-94 ,
-93 ,
-91 ,
-89 ,
-87 ,
-85 ,
-82 ,
-79 ,
-75 ,
-72 ,
-68 ,
-64 ,
-60 ,
-55 ,
-50 ,
-45 ,
-40 ,
-35 ,
-29 ,
-24 ,
-18 ,
-12 ,
-6);

process (CS)
begin
	case CS is	
		when "00" => dataBus <= std_logic_vector(to_signed(to_integer(sine(to_integer(unsigned(address)))), 32));
		when "01" => dataBus <= std_logic_vector(to_signed(to_integer(square(to_integer(unsigned(address)))), 32));
		when "10" => dataBus <= std_logic_vector(to_signed(to_integer(triangle(to_integer(unsigned(address)))), 32));
		when "11" => dataBus <= std_logic_vector(to_signed(to_integer(special(to_integer(unsigned(address)))), 32));
	end case;
end process;
	
end MemArch;	
