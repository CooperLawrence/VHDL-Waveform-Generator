library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity Memory is
port(
	CS: in std_logic_vector(1 downto 0); --Current state
	--EN: in std_logic; --Enable
	address: in std_logic_vector (6 downto 0); -- Address bus
	dataBus: out std_logic_vector(7 downto 0) --Data Bus
	);
end Memory;

architecture MemArch of Memory is
type Sine_array is array (0 to 127) of integer; --look-up table for Sine wave
type Square_array is array (0 to 127) of integer; --look-up table for Square wave
type Triangle_array is array (0 to 127) of integer; --look-up table for Triangle wave
type Special_array is array (0 to 127) of integer; --look-up table for damped-sine wave

signal sine : Sine_array;
signal square : Square_array;
signal triangle : Triangle_array;
signal special : Special_array;



begin
sine <= (0 ,
6 ,
12 ,
18 ,
24 ,
30 ,
36 ,
42 ,
48 ,
54 ,
59 ,
65 ,
70 ,
75 ,
80 ,
85 ,
89 ,
94 ,
98 ,
102 ,
105 ,
108 ,
112 ,
114 ,
117 ,
119 ,
121 ,
123 ,
124 ,
125 ,
126 ,
126 ,
127 ,
126 ,
126 ,
125 ,
124 ,
123 ,
121 ,
119 ,
117 ,
114 ,
112 ,
108 ,
105 ,
102 ,
98 ,
94 ,
89 ,
85 ,
80 ,
75 ,
70 ,
65 ,
59 ,
54 ,
48 ,
42 ,
36 ,
30 ,
24 ,
18 ,
12 ,
6 ,
0 ,
-6 ,
-12 ,
-18 ,
-24 ,
-30 ,
-36 ,
-42 ,
-48 ,
-54 ,
-59 ,
-65 ,
-70 ,
-75 ,
-80 ,
-85 ,
-89 ,
-94 ,
-98 ,
-102 ,
-105 ,
-108 ,
-112 ,
-114 ,
-117 ,
-119 ,
-121 ,
-123 ,
-124 ,
-125 ,
-126 ,
-126 ,
-127 ,
-126 ,
-126 ,
-125 ,
-124 ,
-123 ,
-121 ,
-119 ,
-117 ,
-114 ,
-112 ,
-108 ,
-105 ,
-102 ,
-98 ,
-94 ,
-89 ,
-85 ,
-80 ,
-75 ,
-70 ,
-65 ,
-59 ,
-54 ,
-48 ,
-42 ,
-36 ,
-30 ,
-24 ,
-18 ,
-12 ,
-6);
square <= (127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127 ,
-127);
triangle <= (0 ,
3 ,
7 ,
11 ,
15 ,
19 ,
23 ,
27 ,
31 ,
35 ,
39 ,
43 ,
47 ,
51 ,
55 ,
59 ,
63 ,
67 ,
71 ,
75 ,
79 ,
83 ,
87 ,
91 ,
95 ,
99 ,
103 ,
107 ,
111 ,
115 ,
119 ,
123 ,
127 ,
123 ,
119 ,
115 ,
111 ,
107 ,
103 ,
99 ,
95 ,
91 ,
87 ,
83 ,
79 ,
75 ,
71 ,
67 ,
63 ,
59 ,
55 ,
51 ,
47 ,
43 ,
39 ,
35 ,
31 ,
27 ,
23 ,
19 ,
15 ,
11 ,
7 ,
3 ,
0 ,
-3 ,
-7 ,
-11 ,
-15 ,
-19 ,
-23 ,
-27 ,
-31 ,
-35 ,
-39 ,
-43 ,
-47 ,
-51 ,
-55 ,
-59 ,
-63 ,
-67 ,
-71 ,
-75 ,
-79 ,
-83 ,
-87 ,
-91 ,
-95 ,
-99 ,
-103 ,
-107 ,
-111 ,
-115 ,
-119 ,
-123 ,
0 ,
3 ,
7 ,
11 ,
15 ,
19 ,
23 ,
27 ,
31 ,
35 ,
39 ,
43 ,
47 ,
51 ,
55 ,
59 ,
63 ,
67 ,
71 ,
75 ,
79 ,
83 ,
87 ,
91 ,
95 ,
99 ,
103 ,
107 ,
111 ,
115 ,
119 ,
123);
special <= (0 ,
0 ,
0 ,
0 ,
0 ,
1 ,
1 ,
2 ,
3 ,
3 ,
4 ,
5 ,
6 ,
7 ,
8 ,
9 ,
11 ,
12 ,
13 ,
15 ,
16 ,
17 ,
19 ,
20 ,
21 ,
23 ,
24 ,
25 ,
27 ,
28 ,
29 ,
30 ,
31 ,
32 ,
33 ,
34 ,
35 ,
35 ,
36 ,
36 ,
36 ,
36 ,
36 ,
36 ,
36 ,
35 ,
35 ,
34 ,
33 ,
32 ,
31 ,
30 ,
28 ,
27 ,
25 ,
23 ,
21 ,
19 ,
16 ,
14 ,
11 ,
8 ,
6 ,
3 ,
0 ,
-3 ,
-6 ,
-9 ,
-13 ,
-16 ,
-20 ,
-23 ,
-27 ,
-30 ,
-34 ,
-38 ,
-41 ,
-45 ,
-49 ,
-52 ,
-56 ,
-59 ,
-62 ,
-66 ,
-69 ,
-72 ,
-75 ,
-78 ,
-80 ,
-83 ,
-85 ,
-87 ,
-89 ,
-91 ,
-92 ,
-94 ,
-95 ,
-96 ,
-96 ,
-97 ,
-97 ,
-97 ,
-96 ,
-96 ,
-95 ,
-94 ,
-92 ,
-91 ,
-89 ,
-86 ,
-84 ,
-81 ,
-78 ,
-75 ,
-71 ,
-67 ,
-63 ,
-59 ,
-55 ,
-50 ,
-45 ,
-40 ,
-35 ,
-29 ,
-24 ,
-18 ,
-12 ,
-6);

process (CS)
begin
	case CS is	
		when "00" => dataBus <= std_logic_vector(to_signed(sine(to_integer(unsigned(address))), 8));
		when "01" => dataBus <= std_logic_vector(to_signed(square(to_integer(unsigned(address))), 8));
		when "10" => dataBus <= std_logic_vector(to_signed(triangle(to_integer(unsigned(address))), 8));
		when others => dataBus <= std_logic_vector(to_signed(special(to_integer(unsigned(address))), 8)); -- when "11" gave error of only 4 out of 81 cases covered
	end case;
end process;
	
end MemArch;	
