library ieee;
use ieee.std_logic_1164.all;

entity Memory is
port(
	CS: in std_logic; --Current state?
	EN: in std_logic; --Enable?
	clk: in std_logic; --clock (do we need this?)
	dataBus: out std_logic_vector(31 downto 0); --Data Bus (for the array?)
	address: in std_logic_vector (6 downto 0) -- Address bus
	);
end Memory;

architecture MemArch of Memory is
type Sine_array is array (0 to 127) of float; --look-up table for Sine wave
type Square_array is array (0 to 127) of float; --look-up table for Square wave
type Triangle_array is array (0 to 127) of float; --look-up table for Triangle wave
type Special_array is array (0 to 127) of float; --look-up table for damped-sine wave

begin
Sine_array := (" 0.0 ",
" 0.049067674327418015 ",
" 0.0980171403295606 ",
" 0.14673047445536175 ",
" 0.19509032201612825 ",
" 0.24298017990326387 ",
" 0.29028467725446233 ",
" 0.33688985339222005 ",
" 0.3826834323650898 ",
" 0.4275550934302821 ",
" 0.47139673682599764 ",
" 0.5141027441932217 ",
" 0.5555702330196022 ",
" 0.5956993044924334 ",
" 0.6343932841636455 ",
" 0.6715589548470183 ",
" 0.7071067811865476 ",
" 0.7409511253549591 ",
" 0.7730104533627369 ",
" 0.8032075314806448 ",
" 0.8314696123025452 ",
" 0.8577286100002721 ",
" 0.8819212643483549 ",
" 0.9039892931234433 ",
" 0.9238795325112867 ",
" 0.9415440651830208 ",
" 0.9569403357322089 ",
" 0.970031253194544 ",
" 0.9807852804032304 ",
" 0.989176509964781 ",
" 0.9951847266721968 ",
" 0.9987954562051724 ",
" 1.0 ",
" 0.9987954562051724 ",
" 0.9951847266721969 ",
" 0.989176509964781 ",
" 0.9807852804032304 ",
" 0.970031253194544 ",
" 0.9569403357322089 ",
" 0.9415440651830208 ",
" 0.9238795325112867 ",
" 0.9039892931234434 ",
" 0.881921264348355 ",
" 0.8577286100002721 ",
" 0.8314696123025453 ",
" 0.8032075314806449 ",
" 0.7730104533627371 ",
" 0.740951125354959 ",
" 0.7071067811865476 ",
" 0.6715589548470186 ",
" 0.6343932841636455 ",
" 0.5956993044924335 ",
" 0.5555702330196022 ",
" 0.5141027441932218 ",
" 0.4713967368259978 ",
" 0.42755509343028203 ",
" 0.3826834323650899 ",
" 0.33688985339222033 ",
" 0.2902846772544624 ",
" 0.24298017990326407 ",
" 0.1950903220161286 ",
" 0.1467304744553618 ",
" 0.09801714032956083 ",
" 0.049067674327417966 ",
" 1.2246467991473532e-16 ",
" -0.049067674327417724 ",
" -0.09801714032956059 ",
" -0.14673047445536158 ",
" -0.19509032201612836 ",
" -0.24298017990326382 ",
" -0.2902846772544621 ",
" -0.3368898533922201 ",
" -0.38268343236508967 ",
" -0.4275550934302818 ",
" -0.47139673682599764 ",
" -0.5141027441932216 ",
" -0.555570233019602 ",
" -0.5956993044924332 ",
" -0.6343932841636453 ",
" -0.6715589548470184 ",
" -0.7071067811865475 ",
" -0.7409511253549589 ",
" -0.7730104533627367 ",
" -0.803207531480645 ",
" -0.8314696123025452 ",
" -0.857728610000272 ",
" -0.8819212643483549 ",
" -0.9039892931234431 ",
" -0.9238795325112865 ",
" -0.9415440651830208 ",
" -0.9569403357322088 ",
" -0.970031253194544 ",
" -0.9807852804032303 ",
" -0.9891765099647809 ",
" -0.9951847266721969 ",
" -0.9987954562051724 ",
" -1.0 ",
" -0.9987954562051724 ",
" -0.9951847266721969 ",
" -0.9891765099647809 ",
" -0.9807852804032304 ",
" -0.970031253194544 ",
" -0.9569403357322089 ",
" -0.9415440651830209 ",
" -0.9238795325112866 ",
" -0.9039892931234433 ",
" -0.881921264348355 ",
" -0.8577286100002722 ",
" -0.8314696123025455 ",
" -0.8032075314806453 ",
" -0.7730104533627369 ",
" -0.7409511253549591 ",
" -0.7071067811865477 ",
" -0.6715589548470187 ",
" -0.6343932841636459 ",
" -0.5956993044924332 ",
" -0.5555702330196022 ",
" -0.5141027441932219 ",
" -0.4713967368259979 ",
" -0.42755509343028253 ",
" -0.3826834323650904 ",
" -0.33688985339222 ",
" -0.2902846772544625 ",
" -0.24298017990326418 ",
" -0.19509032201612872 ",
" -0.1467304744553624 ",
" -0.0980171403295605 ",
" -0.04906767432741809 ");
Square_array := (" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" 1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ",
" -1 ");
Triangle_array := ( " 0.0 ",
" 0.03125 ",
" 0.0625 ",
" 0.09375 ",
" 0.125 ",
" 0.15625 ",
" 0.1875 ",
" 0.21875 ",
" 0.25 ",
" 0.28125 ",
" 0.3125 ",
" 0.34375 ",
" 0.375 ",
" 0.40625 ",
" 0.4375 ",
" 0.46875 ",
" 0.5 ",
" 0.53125 ",
" 0.5625 ",
" 0.59375 ",
" 0.625 ",
" 0.65625 ",
" 0.6875 ",
" 0.71875 ",
" 0.75 ",
" 0.78125 ",
" 0.8125 ",
" 0.84375 ",
" 0.875 ",
" 0.90625 ",
" 0.9375 ",
" 0.96875 ",
" 1.0 ",
" 0.96875 ",
" 0.9375 ",
" 0.90625 ",
" 0.875 ",
" 0.84375 ",
" 0.8125 ",
" 0.78125 ",
" 0.75 ",
" 0.71875 ",
" 0.6875 ",
" 0.65625 ",
" 0.625 ",
" 0.59375 ",
" 0.5625 ",
" 0.53125 ",
" 0.5 ",
" 0.46875 ",
" 0.4375 ",
" 0.40625 ",
" 0.375 ",
" 0.34375 ",
" 0.3125 ",
" 0.28125 ",
" 0.25 ",
" 0.21875 ",
" 0.1875 ",
" 0.15625 ",
" 0.125 ",
" 0.09375 ",
" 0.0625 ",
" 0.03125 ",
" 0.0 ",
" -0.03125 ",
" -0.0625 ",
" -0.09375 ",
" -0.125 ",
" -0.15625 ",
" -0.1875 ",
" -0.21875 ",
" -0.25 ",
" -0.28125 ",
" -0.3125 ",
" -0.34375 ",
" -0.375 ",
" -0.40625 ",
" -0.4375 ",
" -0.46875 ",
" -0.5 ",
" -0.53125 ",
" -0.5625 ",
" -0.59375 ",
" -0.625 ",
" -0.65625 ",
" -0.6875 ",
" -0.71875 ",
" -0.75 ",
" -0.78125 ",
" -0.8125 ",
" -0.84375 ",
" -0.875 ",
" -0.90625 ",
" -0.9375 ",
" -0.96875 ",
" 0.0 ",
" 0.03125 ",
" 0.0625 ",
" 0.09375 ",
" 0.125 ",
" 0.15625 ",
" 0.1875 ",
" 0.21875 ",
" 0.25 ",
" 0.28125 ",
" 0.3125 ",
" 0.34375 ",
" 0.375 ",
" 0.40625 ",
" 0.4375 ",
" 0.46875 ",
" 0.5 ",
" 0.53125 ",
" 0.5625 ",
" 0.59375 ",
" 0.625 ",
" 0.65625 ",
" 0.6875 ",
" 0.71875 ",
" 0.75 ",
" 0.78125 ",
" 0.8125 ",
" 0.84375 ",
" 0.875 ",
" 0.90625 ",
" 0.9375 ",
" 0.96875 ");
Special_array := (" 0.0 ",
" 0.00038334120568295324",
" 0.0015315178176493844 ",
" 0.003438995495047541 ",
" 0.006096572563004008 ",
" 0.009491413277471245 ",
" 0.013607094246302923 ",
" 0.018423663857387033 ",
" 0.02391771452281811 ",
" 0.03006246750681671 ",
" 0.03682787006453107 ",
" 0.04418070457910499 ",
" 0.052084709345587704 ",
" 0.06050071061251276 ",
" 0.06938676545539872 ",
" 0.07869831502113496 ",
" 0.08838834764831845 ",
" 0.09840757133620551 ",
" 0.10870459500413487 ",
" 0.11922611795415822 ",
" 0.1299171269222727 ",
" 0.14072110007816965 ",
" 0.1515802173098735 ",
" 0.16243557610811873 ",
" 0.17322741234586625 ",
" 0.18389532523105875 ",
" 0.19437850569560494 ",
" 0.2046159674707241 ",
" 0.21454678008820666 ",
" 0.2241103030388957 ",
" 0.23324642031379614 ",
" 0.2418957745496902 ",
" 0.25 ",
" 0.257501953552896 ",
" 0.2643459430223023 ",
" 0.27047795194349483 ",
" 0.27584586011340856 ",
" 0.28039965912654785 ",
" 0.2840916621704995 ",
" 0.2868767073604517 ",
" 0.2887123539097771 ",
" 0.28955907045360296 ",
" 0.289380414864304 ",
" 0.28814320492196643 ",
" 0.285817679229 ",
" 0.28237764778616425 ",
" 0.2778006316772336 ",
" 0.272067991341274 ",
" 0.26516504294495535 ",
" 0.2570811624023743 ",
" 0.247809876626424 ",
" 0.23734894163370396 ",
" 0.22570040716421338 ",
" 0.21287066751750588 ",
" 0.19887049834846782 ",
" 0.1837150792083243 ",
" 0.16742400165972682 ",
" 0.1500212628387231 ",
" 0.13153524438092826 ",
" 0.11199867667416077 ",
" 0.09144858844506029 ",
" 0.06992624173263336 ",
" 0.047477052347131024 ",
" 0.02415049595802603 ",
" 6.123233995736766e-17 "
" -0.024917178369391814 "
" -0.05054008798242968 ",
" -0.07680423272272832 ",
" -0.10364173357106819 ",
" -0.13098150322910315 ",
" -0.15874943287353396 ",
" -0.18686859055349708 ",
" -0.21525943070536294 ",
" -0.24384001422195759 ",
" -0.2725262384775299 ",
" -0.3012320766757158 ",
" -0.32986982585538865 ",
" -0.3583503628587294 ",
" -0.3865834075372213 ",
" -0.4144777924446442 ",
" -0.44194173824159216 ",
" -0.4688831340136849 ",
" -0.49520982168550315 ",
" -0.5208298836944808 ",
" -0.5456519330735453 ",
" -0.5695854050783057 ",
" -0.592540849484051 ",
" -0.6144302226698403 ",
" -0.6351671786015095 ",
" -0.6546673578225691 ",
" -0.6728486735617093 ",
" -0.6896315940679961 ",
" -0.7049394202898218 ",
" -0.7186985580212861 ",
" -0.7308387836498946 ",
" -0.7412935026522764 ",
" -0.75 ",
" -0.7568996816554822 ",
" -0.7619383063584008 ",
" -0.7650662069258852 ",
" -0.7662385003150238 ",
" -0.7654152857238199 ",
" -0.762561830036604 ",
" -0.7576487399519621 ",
" -0.7506521201654204 ",
" -0.7415537170153246 ",
" -0.7303410470384816 ",
" -0.7170075099221026 ",
" -0.7015524853802727 ",
" -0.683981413526487 ",
" -0.664305858358602 ",
" -0.6425435540187536 ",
" -0.6187184335382292 ",
" -0.5928606398258837 ",
" -0.5650065187082471 ",
" -0.5351985938799205 ",
" -0.5034855236740144 ",
" -0.4699220396141169 ",
" -0.43456886676146683 ",
" -0.3974926259234658 ",
" -0.35876571784227224 ",
" -0.31846618953483297 ",
" -0.2766775830081596 ",
" -0.23348876662579293 ",
" -0.1889937494531247 ",
" -0.14329147896031483 ",
" -0.09648562251191112 ",
" -0.04868433312173514 ");

process (CS)
begin
	case CS is	
		when "00" => dataBus <= Sine_array;
		when "01" => dataBus <= Square_array;
		when "10" => dataBus <= Triangle_array;
		when "11" => dataBus <= Special_array;
	end case;
end process;
	
end MemArch;	
